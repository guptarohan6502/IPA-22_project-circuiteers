module DECODE_REG();

endmodule