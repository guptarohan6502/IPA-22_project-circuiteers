module Processor;






endmodule