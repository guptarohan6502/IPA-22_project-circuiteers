
module split();
endmodule

module Align();
endmodule

module select_PC();
endmodule


