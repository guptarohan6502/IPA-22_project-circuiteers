module Processor;


endmodule