
module PIPE_CONTROL_LOGIC();





endmodule