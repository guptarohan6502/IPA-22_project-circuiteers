module FETCH_REG(predict_pc, F_pred_PC);


endmodule


